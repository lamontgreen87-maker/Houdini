// Gatling V1: AXI-Lite Wrapper for 16-Channel Matrix Capture
// Maps the 4x4 Grid results to the Zynq Memory Map

module gatling_axi_wrapper # (
    parameter integer C_S_AXI_DATA_WIDTH = 32,
    parameter integer C_S_AXI_ADDR_WIDTH = 7   // Enough space for 16 channels + control
)(
    // AXI-Lite Interface Signals
    input  wire  S_AXI_ACLK,
    input  wire  S_AXI_ARESETN,
    input  wire [C_S_AXI_ADDR_WIDTH-1 : 0] S_AXI_AWADDR,
    input  wire  S_AXI_AWVALID,
    output wire  S_AXI_AWREADY,
    input  wire [C_S_AXI_DATA_WIDTH-1 : 0] S_AXI_WDATA,
    input  wire  S_AXI_WVALID,
    output wire  S_AXI_WREADY,
    output wire [1 : 0] S_AXI_BRESP,
    output wire  S_AXI_BVALID,
    input  wire  S_AXI_BREADY,
    input  wire [C_S_AXI_ADDR_WIDTH-1 : 0] S_AXI_ARADDR,
    input  wire  S_AXI_ARVALID,
    output wire  S_AXI_ARREADY,
    output wire [C_S_AXI_DATA_WIDTH-1 : 0] S_AXI_RDATA,
    output wire [1 : 0] S_AXI_RRESP,
    output wire  S_AXI_RVALID,
    input  wire  S_AXI_RREADY,

    // External Connections to the Sensors
    input  wire [15:0] adc_raw_in,
    input  wire        adc_sync
);

    // Instantiate the Capture Engine we drafted earlier
    wire [11:0] channel_out [0:15];
    wire data_ready;
    reg trigger;

    adc_capture_engine engine_inst (
        .clk(S_AXI_ACLK),
        .reset_n(S_AXI_ARESETN),
        .adc_data_in(adc_raw_in),
        .adc_frame_sync(adc_sync),
        .trigger_capture(trigger),
        .channel_buffer(channel_out),
        .data_valid(data_ready)
    );

    // --- AXI Read Logic ---
    // This allows Python to "see" the 16 channels as registers 0-15
    assign S_AXI_RDATA = (S_AXI_ARADDR[5:2] < 16) ? channel_out[S_AXI_ARADDR[5:2]] : 32'hDEADBEEF;

    // --- AXI Write Logic ---
    // Writing to register 16 toggles the trigger
    always @(posedge S_AXI_ACLK) begin
        if (S_AXI_WVALID && S_AXI_AWADDR[6:2] == 16) 
            trigger <= S_AXI_WDATA[0];
        else 
            trigger <= 0;
    end

    // (Simplified AXI handshake logic below - usually generated by Vivado IP Integrator)
    assign S_AXI_AWREADY = 1'b1;
    assign S_AXI_WREADY  = 1'b1;
    assign S_AXI_ARREADY = 1'b1;
    assign S_AXI_RVALID  = 1'b1;
    assign S_AXI_BVALID  = 1'b1;

endmodule
